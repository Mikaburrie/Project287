module Project287(input a, output reg b);

	always @(*) begin
	
		b = a;
	
	end

endmodule
