module counter_inc1();

	

endmodule
